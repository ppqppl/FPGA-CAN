module can_top(
    input   wire    clk     ,
    input   wire    rstn    ,

    input   wire    can_h   ,
    input   wire    can_l

);



endmodule